module DecToBin(D9, D8, D7, D6, D5, D4, D3, D2, D1, D0, Y4, Y3, Y2, Y0);

input D9, D8, D7, D6, D5, D4, D3, D2, D1, D0;
output reg Y4, Y3, Y2, Y0;

always @(*) begin
    
    case ({D9, D8, D7, D6, D5, D4, D3, D2, D1, D0})
        10'b00_0000_0001: {Y4, Y3, Y2, Y0} = 4'b0000; 
        10'b00_0000_0010: {Y4, Y3, Y2, Y0} = 4'b0001;
        10'b00_0000_0100: {Y4, Y3, Y2, Y0} = 4'b0010;
        10'b00_0000_1000: {Y4, Y3, Y2, Y0} = 4'b0011;
        10'b00_0001_0000: {Y4, Y3, Y2, Y0} = 4'b0100;
        10'b00_0010_0000: {Y4, Y3, Y2, Y0} = 4'b0101;
        10'b00_0100_0000: {Y4, Y3, Y2, Y0} = 4'b0110;
        10'b00_1000_0000: {Y4, Y3, Y2, Y0} = 4'b0111;
        10'b01_0000_0000: {Y4, Y3, Y2, Y0} = 4'b1000;
        10'b10_0000_0000: {Y4, Y3, Y2, Y0} = 4'b1001;
        default: {Y4, Y3, Y2, Y0} = 4'd0;
    endcase

end

endmodule